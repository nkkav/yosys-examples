module and2(f, a, b);
  output f;
  input a, b;
  
  assign f = a & b;

endmodule
